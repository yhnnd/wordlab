<#gry-#gry>(
<#gry-#gry>( )<-wte>(name = "inanimate objects"
<#gry-#gry>( )<-wte>(value = "things that are not alive"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
