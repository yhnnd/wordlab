<-wte>(function system <"main"><blu-wte>(go back);
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
