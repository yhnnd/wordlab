<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "multimedia data objects"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
