<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "a noun or pronoun representing the person or thing that something is done to"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
