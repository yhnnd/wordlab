<-wte>(<"object-word"><-ylw>(word                                          )
<-wte>(
<-wte>(<"object-sort[1]"><-ylw>(sort[1]                                       )  <"object-sort[1].def[1]"><-ylw>(sort[1].def[1]                                )
<-wte>(<"object-sort[1].def[1].example[1]"><-ylw>(sort[1].def[1].example[1]                     )  <"object-sort[1].def[1].example[2]"><-ylw>(sort[1].def[1].example[2]                     )
<-wte>(<"object-sort[1].def[1].example[3]"><-ylw>(sort[1].def[1].example[3]                     )  <"object-sort[1].def[1].example[3].explaination[1]"><-ylw>(sort[1].def[1].example[3].explaination[1]     )
<-wte>(<"object-sort[1].def[2]"><-ylw>(sort[1].def[2]                                )  <"object-sort[1].def[2].also[1]"><-ylw>(sort[1].def[2].also[1]                        )
<-wte>(<"object-sort[1].def[2].also[2]"><-ylw>(sort[1].def[2].also[2]                        )  <"object-sort[1].def[2].example[1]"><-ylw>(sort[1].def[2].example[1]                     )
<-wte>(<"object-sort[1].def[2].example[2]"><-ylw>(sort[1].def[2].example[2]                     )  <"object-sort[1].def[2].example[3]"><-ylw>(sort[1].def[2].example[3]                     )
<-wte>(<"object-sort[1].def[2].example[3].explaination[1]"><-ylw>(sort[1].def[2].example[3].explaination[1]     )  <"object-sort[1].def[3]"><-ylw>(sort[1].def[3]                                )
<-wte>(<"object-sort[1].def[3].also[1]"><-ylw>(sort[1].def[3].also[1]                        )  <"object-sort[1].def[4]"><-ylw>(sort[1].def[4]                                )
<-wte>(<"object-sort[1].def[4].example[1]"><-ylw>(sort[1].def[4].example[1]                     )  
<-wte>(
<-wte>(<"object-sort[2]"><-ylw>(sort[2]                                       )  <"object-sort[2].def[1]"><-ylw>(sort[2].def[1]                                )
<-wte>(<"object-sort[2].def[1].example[1]"><-ylw>(sort[2].def[1].example[1]                     )  <"object-sort[2].def[1].example[2]"><-ylw>(sort[2].def[1].example[2]                     )
<-wte>(<"object-sort[2].def[1].example[3]"><-ylw>(sort[2].def[1].example[3]                     )  
<-wte>(
<-wte>(<"object-sort[3]"><-ylw>(sort[3]                                       )  <"object-sort[3].def[1]"><-ylw>(sort[3].def[1]                                )
<-wte>(<"object-sort[3].def[1].example[1]"><-ylw>(sort[3].def[1].example[1]                     )  <"object-sort[3].def[1].example[2]"><-ylw>(sort[3].def[1].example[2]                     )
<-wte>(<blu-blu>(
