<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "If no one objects, I would like Mrs Harrison to be present."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
