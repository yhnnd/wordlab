<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "the purpose of a plan, action, or activity"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
