<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "an everyday object such as a spoon"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
