Search;
<-gry>(cannot locate) <-ylw>(database damaged line);
<-gry>(cannot translate) <-ylw>(redirected words);
<-gry>(cannot record) <-ylw>(translating history);
<-gry>(cannot record) <-ylw>(translating error);
<-gry>(cannot support) <-ylw>(translating rules);
<-gry>(cannot add) <-red>(affixes) <-cyn>(special words) <-grn>(rules);
<-ylw>(WOC1 do for)<-gry>(error placing) <-ylw>(do) <-gry>(when nothing after) <-ylw>(for);
<-ylw>(Word Cutter)<-gry>(cannot translate words with) <-ylw>(multiple affixes);



