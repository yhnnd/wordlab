<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "n."
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
