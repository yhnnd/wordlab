<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "to play a trump that beats someone else's card in a game"                            <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "出王牌赢\(在游戏中打出击败别人的牌的王牌\);"                        <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
