<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "goal"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
