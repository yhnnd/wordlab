<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "to play a trump that beats someone else's card in a game"
<#gry-#gry>( )<-wte>(Chinese = "[�����[����]��������A[�e�˵���];"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
