<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "object"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
