<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "v."                                                                                    <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
