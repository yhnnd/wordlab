<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "trump"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
