<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "a noun or pronoun representing the person or thing that something is done to"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
