<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "a small metal object"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
