<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "vt."
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
