<-wte>(const char *cmd_funct[]
<-gry>("cmd_funct:","select","create","delete","insert","update","fetch","drop","add"
<-gry>("open","set","alter","order_by","group_by","print","system","join","check","#"
<-wte>(const char *cmd_scope[]
<-gry>("cmd_scope:","where","from","to","in","between","of","#"
<-wte>(const char *cmd_conj []
<-gry>("cmd_conj:","and","or","not","if","else","#"
<-wte>(const char *cmd_data []
<-gry>("cmd_data:","library","source","#"
<-wte>(<"main"><blu-wte>(go back)
