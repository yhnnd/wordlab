<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "��My name��s not Sonny,�� the child objected."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
