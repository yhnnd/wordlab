<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "Robson strongly objected to the terms of the contract."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
