 Do you mean apply ?
 Do you mean apply ?
 Do you mean apply ?
<red-> (error) <ylw->(\(illegal choice\))
 Do you mean apply ?
 Do you mean apply ?
 Do you mean apply ?
 Do you mean apply ?
 Do you mean apply ?
press [A] to add <fore yellow>(qqfsdf
)
press [D] to delete <fore red>(qqfsdf
)
press [U] to update <fore cyan>(qqfsdf
)
