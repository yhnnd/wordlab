<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "By wearing a simple but stunning dress, she had trumped them all."
<#gry-#gry>( )<-wte>(Chinese = "������һ�l���΅s�@�G��ȹ��,����Ⱥ��."
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
