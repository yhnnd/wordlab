<blk-gry>(<#red-gry>(Add Word Files/Settings/WL/addword                         );
<blk-wte>(<button="setWord"><-wte>(word)<gry-wte>( word to add)<-wte>(                                           );
<blk-gry>(<#red-gry>(Add Definition                                             );
<blk-wte>(<button="setSort"><-wte>(sort)<gry-wte>( $def_sort)<-wte>(                                             );
<blk-gry>(<button="setTrans"><-wte>(definition)<gry-wte>( $def_trans)<-wte>(                                      );
<blk-wte>(<button="addDef"><-ylw>( add definition  )<button="resetDef"><ylw-red>( reset definition )<gry-wte>(                        );
<blk-gry>(<#red-gry>(Save All Definitions                                       );
<blk-wte>(<button="addAllDefs"><-ylw>( add all defintions  )<button="resetAllDefs"><ylw-red>( reset all definitions )<gry-wte>(               );
<blk-gry>(<button="printAllDefs"><gry-wte>( print all defs )<gry-wte>( $defs                                     );
<blk-wte>(<button="printAllData"><-cyn>( print all data )<#blu-wte>( developed by skyside inc. 2016/12/09      );
