<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "to state a fact or opinion as a reason for opposing or disapproving of something"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
