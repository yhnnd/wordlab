<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "My object was to explain the decision simply."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
