<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "If no one objects, I would like Mrs Harrison to be present."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
