<#blu-#blu>(
<#blu-#blu>( )<-wte>(name = "suit"                                                                                   <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(value = "one of the four types of cards in a set"                                               <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
