<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "to state a fact or opinion as a reason for opposing or disapproving of something"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
