<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "object"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
