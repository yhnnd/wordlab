<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "But then he decided to play his trump card."                                         <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "但后来他决定打出自己的王牌."                                            <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
