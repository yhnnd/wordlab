<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "scientists studying plants, animals, or inanimate objects"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
