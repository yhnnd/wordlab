<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "The object of the game is to improve children��s math skills."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
