<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "I objected to having to rewrite the article."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
