<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "a combination of written information on a computer and instructions that act on the inf
<#gry-#gry>( )<-wte>(ormation, for example in the form of a document or a picture"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
