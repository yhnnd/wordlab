<#blu-#blu>(
<#blu-#blu>( )<-wte>(name = "the object of the exercise"
<#blu-#blu>( )<-wte>(value = "the purpose of what you are doing"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
