<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "the suit chosen to have a higher value than the other suits in a particular card game"
<#gry-#gry>( )<-wte>(Chinese = "[�����[���е�]���ƻ�ɫ;"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
