<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "direct object"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
