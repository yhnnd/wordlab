<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "The group objected that the policy would prevent patients from receiving the best treat
<#blu-#blu>( )<-wte>(ment."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
