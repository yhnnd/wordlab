<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "trumps"                                                                                <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
