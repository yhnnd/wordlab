<#blu-#blu>(
<#blu-#blu>( )<-wte>(name = "play his trump card"                                                                    <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(value = "use his advantage"                                                                     <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
