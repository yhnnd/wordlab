<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "aim"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
