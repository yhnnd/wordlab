<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "to feel or say that you oppose or disapprove of something"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
