<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "vi."
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
