<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "scientists studying plants, animals, or inanimate objects"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
