<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "to do better than someone else in a situation when people are competing with each oth<#blu-#blu>(  )
<#blu-#blu>( )<-wte>(er"                                                                                             <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "胜过;打败;发挥出色;掌握主动权;"                                         <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
