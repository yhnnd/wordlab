<#gry-#gry>(
<#gry-#gry>( )<-wte>(name = "They hold all the trump cards"
<#gry-#gry>( )<-wte>(value = "They have things which could give them an advantage"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
