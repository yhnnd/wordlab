<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "Hearts are the trumps."                                                              <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "红桃是王牌."                                                                    <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
