<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "n."
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
