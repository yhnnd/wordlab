<-wte>(
<-gry>(
<-gry>(
<-wte>(
<-gry>(
<-gry>(
<-wte>(
<-gry>(
<-gry>(
<-wte>(<"system info"><blu-wte>(go back)
