<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "trump"                                                                                 <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
