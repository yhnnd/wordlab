<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "I objected to having to rewrite the article."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
