<#gry-#gry>(
<#gry-#gry>( )<-wte>(name = "the object of the exercise"
<#gry-#gry>( )<-wte>(value = "the purpose of what you are doing"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
