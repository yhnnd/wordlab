<#gry-#gry>(
<#gry-#gry>( )<-wte>(name = "suit"
<#gry-#gry>( )<-wte>(value = "one of the four types of cards in a set"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
