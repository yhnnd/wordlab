<blk-gry>(<#red-gry>(Add Word) <#blu-gry>(Files/Settings/WL/addword;
<blk-wte>(<button="setWord"><-wte>(word)<gry-wte>( $word )<-wte>(;
<blk-gry>(<#red-gry>(Add Definition;
<blk-wte>(<button="setSort"><-wte>(sort)<gry-wte>( $def_sort )<-wte>(;
<blk-gry>(<button="setTrans"><-wte>(definition)<gry-wte>( $def_trans )<-wte>(;
<blk-wte>(<button="addDef"><-ylw>( add definition  )<button="resetDef"><ylw-red>( clear )<gry-wte>(;
<blk-gry>(<-gry>(definitions)<wte-gry>( $defs_buf )<-gry>(;
<blk-wte>(<#red-gry>(Save All Definitions;
<blk-gry>(<button="addAllDefs"><-ylw>( Save all defintions  )<button="resetAllDefs"><ylw-red>( delete saved definitions )<gry-wte>(;
<blk-wte>(<button="printAllDefs"><gry-wte>( print all defs )<gry-wte>( $defs_out )<gry-wte>(;
<blk-gry>(<button="printAllData"><-cyn>( print all data );
<blk-wte>(<button="printAllScriptLines"><-cyn>( print all scripts )<#blu-gry>( developed by skyside inc. 2016/12/09;
;