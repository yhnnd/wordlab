<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "to feel or say that you oppose or disapprove of something"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
