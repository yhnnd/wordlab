<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "vt."
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
