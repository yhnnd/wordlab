<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "a solid thing that you can hold, touch, or see but that is not alive"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
