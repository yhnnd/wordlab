<-wte>(
<-gry>(
<-gry>(
<-wte>(
<-gry>(
<-gry>(
<-wte>(
<-gry>(
<-gry>(
<-wte>(<"main"><blu-wte>(go back)
