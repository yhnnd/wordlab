<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "They hold all the trump cards."                                                      <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "他们掌握着所有的王牌."                                                     <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
