<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "to do better than someone else in a situation when people are competing with each other
<#gry-#gry>( )<-wte>("
<#gry-#gry>( )<-wte>(Chinese = "�A;���^;��;"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
