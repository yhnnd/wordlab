<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "By wearing a simple but stunning dress, she had trumped them all."                   <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "通过穿着简单但令人惊叹的衣服,她胜过了所有人."                   <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
