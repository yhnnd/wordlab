<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "a card from the suit that has been chosen to have a higher value than the other suits i
<#gry-#gry>( )<-wte>(n a particular card game"
<#gry-#gry>( )<-wte>(Chinese = "����;����;"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
