<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "vi."
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
