<-wte>(<button="test_print_all_data"><-wte>(show all data);
<-wte>(<button="InitArrayByDeclaration"><-wte>(init array);
<-wte>(<button="InitArrayByLoop1"><-wte>(init array loop 1);
<-wte>(<button="InitArrayByLoop2"><-wte>(init array loop 2);
<-wte>(<button="CreateClass"><-wte>(create class);
;
;
;
;
<-wte>(skyside tech inc.);
#date 2017.03.20.02:51
done;