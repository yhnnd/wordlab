<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "an everyday object such as a spoon"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
