<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "the purpose of a plan, action, or activity"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
