<-wte>(function select <"main"><blu-wte>(go back);
<wte-gry>(;
<-wte>(from/to;
<wte-gry>(select from lth=3 to lth=4;
<-wte>(where name=value;
<wte-gry>(select where sort=n.;
<-wte>(where name=value more;
<wte-gry>(select where index=emp begin=esp end=sion;
<-wte>(in/of;
<wte-gry>(select in word:en-ch;
