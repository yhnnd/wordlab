<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "But then he decided to play his trump card."
<#gry-#gry>( )<-wte>(Chinese = "���^���Q��ʹ�����Ě����."
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
