<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "Robson strongly objected to the terms of the contract."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
