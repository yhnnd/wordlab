<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "a combination of written information on a computer and instructions that act on the inf
<#blu-#blu>( )<-wte>(ormation, for example in the form of a document or a picture"
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
