<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "a small metal object"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
