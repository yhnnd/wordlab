<-wte>(<"trump-word"><-ylw>(word                                          )
<-wte>(
<-wte>(<"trump-sort[1]"><-ylw>(sort[1]                                       )  <"trump-sort[1].def[1]"><-ylw>(sort[1].def[1]                                )
<-wte>(<"trump-sort[1].def[1].explaination[1]"><-ylw>(sort[1].def[1].explaination[1]                )  <"trump-sort[1].def[1].also[1]"><-ylw>(sort[1].def[1].also[1]                        )
<-wte>(<"trump-sort[1].def[1].example[1]"><-ylw>(sort[1].def[1].example[1]                     )  <"trump-sort[1].def[2]"><-ylw>(sort[1].def[2]                                )
<-wte>(<"trump-sort[1].def[2].explaination[1]"><-ylw>(sort[1].def[2].explaination[1]                )  <"trump-sort[1].def[2].also[1]"><-ylw>(sort[1].def[2].also[1]                        )
<-wte>(<"trump-sort[1].def[3]"><-ylw>(sort[1].def[3]                                )  <"trump-sort[1].def[3].also[1]"><-ylw>(sort[1].def[3].also[1]                        )
<-wte>(<"trump-sort[1].def[3].example[1]"><-ylw>(sort[1].def[3].example[1]                     )  <"trump-sort[1].def[3].example[1].explaination[1]"><-ylw>(sort[1].def[3].example[1].explaination[1]     )
<-wte>(<"trump-sort[1].def[3].example[2]"><-ylw>(sort[1].def[3].example[2]                     )  <"trump-sort[1].def[3].example[2].explaination[1]"><-ylw>(sort[1].def[3].example[2].explaination[1]     )
<-wte>(
<-wte>(<"trump-sort[2]"><-ylw>(sort[2]                                       )  <"trump-sort[2].def[1]"><-ylw>(sort[2].def[1]                                )
<-wte>(<"trump-sort[2].def[2]"><-ylw>(sort[2].def[2]                                )  <"trump-sort[2].def[2].example[1]"><-ylw>(sort[2].def[2].example[1]                     )
<-wte>(<blu-blu>(
