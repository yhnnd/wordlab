<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "v."
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
