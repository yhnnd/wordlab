<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "n."                                                                                    <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
