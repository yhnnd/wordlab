<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "trumps"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
