<#blu-#blu>(
<#blu-#blu>( )<-wte>(name = "inanimate objects"
<#blu-#blu>( )<-wte>(value = "things that are not alive"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
