<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "Hearts are the trumps."
<#gry-#gry>( )<-wte>(Chinese = "�t��������"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
