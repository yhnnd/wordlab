<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "trump card"                                                                            <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
