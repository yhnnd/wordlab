<-wte>(function system <"system info"><blu-wte>(go back);
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
<-wte>(;
<-gry>(;
