<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "multimedia data objects"
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
