<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "the suit chosen to have a higher value than the other suits in a particular card game<#blu-#blu>(  )
<#blu-#blu>( )<-wte>("                                                                                               <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "王牌\(花色\);將牌\(花色\);"                                                      <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
