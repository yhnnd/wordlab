<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "direct object"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
