<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "a solid thing that you can hold, touch, or see but that is not alive"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
