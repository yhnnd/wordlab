<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "a card from the suit that has been chosen to have a higher value than the other suits<#blu-#blu>(  )
<#blu-#blu>( )<-wte>( in a particular card game"                                                                     <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(Chinese = "王牌;將牌;"                                                                      <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
