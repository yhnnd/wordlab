<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "The object of the game is to improve children��s math skills."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
