<#blu-#blu>(
<#blu-#blu>( )<-wte>(name = "They hold all the trump cards"                                                          <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(value = "They have things which could give them an advantage"                                   <#blu-#blu>(  )
<#blu-#blu>( )<-wte>(<"trump-main"><-ylw>( go back )
<#blu-#blu>(
