<#gry-#gry>(
<#gry-#gry>( )<-wte>(name = "play his trump card"
<#gry-#gry>( )<-wte>(value = "use his advantage"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
