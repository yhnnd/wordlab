<#blu-#blu>(
<#blu-#blu>( )<-wte>(English = "My object was to explain the decision simply."
<#blu-#blu>( )<-wte>(Chinese = ""
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
