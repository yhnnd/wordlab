<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "The customer will benefit most, and that is the object of the exercise."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
