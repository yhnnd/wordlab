<#gry-#gry>(
<#gry-#gry>( )<-wte>(English = "The group objected that the policy would prevent patients from receiving the best treat
<#gry-#gry>( )<-wte>(ment."
<#gry-#gry>( )<-wte>(Chinese = ""
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
