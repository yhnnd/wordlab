<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "aim"
<#gry-#gry>( )<-wte>(<"object-main"><-ylw>( go back )
<#gry-#gry>(
