<#blu-#blu>(
<#blu-#blu>( )<-wte>(value = "goal"
<#blu-#blu>( )<-wte>(<"object-main"><-ylw>( go back )
<#blu-#blu>(
