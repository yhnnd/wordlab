<#gry-#gry>(
<#gry-#gry>( )<-wte>(value = "trump card"
<#gry-#gry>( )<-wte>(<"trump-main"><-ylw>( go back )
<#gry-#gry>(
